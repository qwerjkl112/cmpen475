`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/12/2017 04:43:09 PM
// Design Name: 
// Module Name: carry_look_ahead
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: x
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module carry_look_ahead128(
input [127:0] a, b,
input clk, cin, 
output [127:0] s, 
output cout    
    );
    
wire c16, c32, c48, c64, c80, c96, c112, ccout;
reg [127:0] rega, regb;

always @ (posedge clk) begin
    rega <= a;
    regb <= b;
end

    	claadder16 m1(rega[15:0], regb[15:0], cin, s[15:0], c16);
        claadder16 m2(rega[31:16], regb[31:16], c16, s[31:16], c32);
        claadder16 m3(rega[47:32], regb[47:32], c32, s[47:32], c48);
        claadder16 m4(rega[63:48], regb[63:48], c48, s[63:48], c64);
        claadder16 m5(rega[79:64], regb[79:64], c64, s[79:64], c80);
        claadder16 m6(rega[95:80], regb[95:80], c80, s[95:80], c96);
        claadder16 m7(rega[111:96], regb[111:96], c96, s[111:96], c112);
        claadder16 m8(rega[127:112], regb[127:112], c112, s[127:112], cout);
endmodule


module claadder16(
input [15:0] a, b,
input cin,
output [15:0] s, 
output cout);

reg tempa, tempb;
wire c1, c2, c3;


claadder4 cla1(a[3:0], b[3:0], cin, s[3:0], c1);
claadder4 cla2(a[7:4], b[7:4], c1, s[7:4], c2);
claadder4 cla3(a[11:8], b[11:8], c2, s[11:8], c3);
claadder4 cla4(a[15:12], b[15:12], c3, s[15:12], cout);

endmodule

module claadder4(
input [3:0] a, b,
input cin,
output [3:0] s, 
output cout);

wire c1, c2, c3, c4, p1, p2, p3, p4, g1, g2, g3, g4;


   assign g1 = a[0] & b[0];
   assign p1 = a[0] | b[0];
   assign g2 = a[1] & b[1];
   assign p2 = a[1] | b[1];   
   assign g3 = a[2] & b[2];
   assign p3 = a[2] | b[2];
   assign g4 = a[3] & b[3];
   assign p4 = a[3] | b[3];
   
   assign c1 = g1 | (p1 & cin);
   assign c2 = g2 | (p2 & g1) | (p2 & p1 & cin);
   assign c3 = g3 | (p3 & g2) | (p3 & p2 & g1) | (p3 & p2 & p1 & cin);
   assign c4 = g4 | (p4 & g3) | (p4 & p3 & g2) | (p4 & p3 & p2 & g1) | (p4 & p3 & p2 & p1 & cin);
   assign cout = c4;
      
   assign s[0] = g1 ^ p1 ^ cin;
   assign s[1] = g2 ^ p2 ^ c1;
   assign s[2] = g3 ^ p3 ^ c2;
   assign s[3] = g4 ^ p4 ^ c3;
   
endmodule
